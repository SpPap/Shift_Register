--Implementation of shift register 24-bit using 6 shift registers 4-bit
--Structural modeling

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY SHIFT_REG24 IS
    
    PORT (
        D : IN STD_LOGIC_VECTOR(0 TO 23); --PARALLEL LOAD
        S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        MR : IN STD_LOGIC; --MASTER RESET (ACTIVE LOW)
        CP : IN STD_LOGIC; --CLOCK
        DSL, DSR : IN STD_LOGIC; --SHIFT LEFT/RIGHT
        Q : BUFFER STD_LOGIC_VECTOR(0 TO 23) --OUTPUT
    );

END ENTITY;

ARCHITECTURE S1 OF SHIFT_REG24 IS

    COMPONENT SHIFT_REG4 IS
        PORT (
            D : IN STD_LOGIC_VECTOR(0 TO 3); --PARALLEL LOAD
            S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
            MR : IN STD_LOGIC; --MASTER RESET (ACTIVE LOW)
            CP : IN STD_LOGIC; --CLOCK
            DSL, DSR : IN STD_LOGIC; --SHIFT LEFT/RIGHT
            Q : BUFFER STD_LOGIC_VECTOR(0 TO 3) --OUTPUT
        );
    END COMPONENT;
	 
	 SIGNAL R0Q : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R1Q : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R2Q : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R3Q : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R4Q : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R5Q : STD_LOGIC_VECTOR(0 TO 3);
	  
	 SIGNAL R0D : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R1D : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R2D : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R3D : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R4D : STD_LOGIC_VECTOR(0 TO 3);
	 SIGNAL R5D : STD_LOGIC_VECTOR(0 TO 3);
	 
    BEGIN
    R0: SHIFT_REG4 PORT MAP(R0D, S, MR, CP, R1Q(0), DSR, R0Q);
    R1: SHIFT_REG4 PORT MAP(R1D, S, MR, CP, R2Q(0),  R0Q(3), R1Q);
    R2: SHIFT_REG4 PORT MAP(R2D, S, MR, CP, R3Q(0), R1Q(3), R2Q);
    R3: SHIFT_REG4 PORT MAP(R3D, S, MR, CP, R4Q(0), R2Q(3), R3Q);
    R4: SHIFT_REG4 PORT MAP(R4D, S, MR, CP, R5Q(0), R3Q(3), R4Q);
    R5: SHIFT_REG4 PORT MAP(R5D, S, MR, CP, DSL, R4Q(3), R5Q);
   
	 
	 Q <= R0Q & R1Q & R2Q & R3Q & R4Q & R5Q; --routing
	

END ARCHITECTURE;